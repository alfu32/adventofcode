module main

pub
