module main

import arrays

fn test_scd(){

	test_cards := "
		Card 1: 41 48 83 86 17 | 83 86  6 31 17  9 48 53
		Card 2: 13 32 20 16 61 | 61 30 68 82 17 32 24 19
		Card 3:  1 21 53 59 44 | 69 82 63 72 16 21 14  1
		Card 4: 41 92 73 84 69 | 59 84 76 51 58  5 54 83
		Card 5: 87 83 26 28 32 | 88 30 70 12 93 22 82 36
		Card 6: 31 18 13 56 72 | 74 77 10 23 35 67 36 11
	".trim_indent()
	println(test_cards)

	cards := test_cards.split("\n").map(card_from_string(it))
	println(cards)
	points := cards.map(it.points())
	println(points)

	mut copies := arrays.flat_map()(cards, fn[cards](c Card) []Card {
		times:=c.points()
		if times > 0 {
			i := c.number
			mut k:=i
			for _ in 1..(times+1) {
				if k >=cards.len {
					k=i
				}
				ctc := arrays.filter(cards,fn [c](c0 Card) bool {
					return c0.number == c.number
				}).map(fn(cc Card) Card {
					Card{
						number: c.number
						code: c.code
						winning_numbers: cc.winning_numbers
						chosen_numbers: cc.chosen_numbers
					}
				})
				k++
				return ctc
			}
		}
	})

}
